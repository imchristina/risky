module risky_writeback (
  input clk,
  output [4:0] reg_sel,
  output [31:0] reg_data
);

endmodule
