// TODO all of this, makefile integration, etc

module risky_tests ();
  // Run all tests

endmodule

module risky_tests_alu ();

endmodule
