module risky_mem (
  input clk
);

endmodule
